Quarter,Time,Down,ToGo,Location,NYG,ATL,Detail,EPB,EPA
,,,,,,,Giants won the coin toss and deferred Falcons to receive the opening kickoff.,,
1,15:00,,,NYG 35,0,0,Graham Gano kicks off 65 yards touchback.,0.000,0.940
1,15:00,1,10,ATL 30,0,0,Michael Penix pass incomplete short left intended for Ray-Ray McCloud (defended by Deonte Banks),0.940,0.390
1,14:52,2,10,ATL 30,0,0,Bijan Robinson right tackle for 3 yards (tackle by Micah McFadden),0.390,0.100
1,14:14,3,7,ATL 33,0,0,Michael Penix pass complete short middle to Drake London for 19 yards (tackle by Adoree' Jackson and Jason Pinnock),0.100,2.390
1,13:33,1,10,NYG 48,0,0,Penalty on Brian Burns: Neutral Zone Infraction 5 yards (accepted) (no play),2.390,3.120
1,13:18,1,5,NYG 43,0,0,Bijan Robinson left tackle for 10 yards (tackle by Darius Muasau),3.120,3.380
1,12:38,1,10,NYG 33,0,0,Michael Penix pass incomplete short left intended for Drake London,3.380,2.840
1,12:34,2,10,NYG 33,0,0,Ray-Ray McCloud right end for 8 yards (tackle by Darius Muasau and Jason Pinnock),2.840,3.200
1,11:52,3,2,NYG 25,0,0,Michael Penix pass incomplete deep right intended for Drake London,3.200,1.930
1,11:48,4,2,NYG 25,0,0,Riley Patterson 43 yard field goal no good,1.930,-1.140
1,11:44,1,10,NYG 33,0,0,Drew Lock pass complete short right to Malik Nabers for 6 yards (tackle by Mike Hughes and Kaden Elliss),1.140,1.400
1,11:05,2,4,NYG 39,0,0,Drew Lock pass incomplete short right,1.400,0.700
1,10:57,3,4,NYG 39,0,0,Drew Lock pass incomplete short right intended for Wan'Dale Robinson,0.700,-0.780
1,10:52,4,4,NYG 39,0,0,Jamie Gillan punts 51 yards fair catch by Avery Williams at ATL-10,-0.780,0.380
1,10:45,1,10,ATL 10,0,0,Bijan Robinson right tackle for 7 yards (tackle by Elijah Chatman),-0.380,-0.090
1,10:08,2,3,ATL 17,0,0,Bijan Robinson left end for 7 yards (tackle by Andru Phillips),-0.090,0.540
1,9:41,1,10,ATL 24,0,0,Michael Penix pass incomplete short right intended for Charlie Woerner,0.540,0.000
1,9:38,2,10,ATL 24,0,0,Michael Penix pass complete short left to Drake London for 5 yards (tackle by Dane Belton and Darius Muasau),0.000,-0.030
1,8:56,3,5,ATL 29,0,0,Michael Penix scrambles right guard for 1 yard (tackle by Kayvon Thibodeaux),-0.030,-1.370
1,8:15,4,4,ATL 30,0,0,Bradley Pinion punts 46 yards returned by Ihmir Smith-Marsette for 6 yards (tackle by Natrone Brooks),-1.370,-0.940
1,8:05,1,10,NYG 30,0,0,Tyrone Tracy right tackle for 4 yards (tackle by David Onyemata),0.940,0.930
1,7:29,2,6,NYG 34,0,0,Drew Lock pass complete short left to Malik Nabers for 6 yards (tackle by Kaden Elliss and Demone Harris),0.930,1.600
1,6:57,1,10,NYG 40,0,0,Drew Lock pass complete short left to Tyrone Tracy for 9 yards (tackle by Justin Simmons),1.600,2.270
1,6:18,2,1,NYG 49,0,0,Tyrone Tracy right tackle for 5 yards (tackle by David Onyemata and Grady Jarrett),2.270,2.520
1,5:34,1,10,ATL 46,0,0,Devin Singletary right tackle for 5 yards (tackle by AJ Terrell and Kaden Elliss),2.520,2.650
1,4:55,2,5,ATL 41,0,0,Devin Singletary left tackle for 4 yards (tackle by Kentavius Street),2.650,2.480
1,4:19,3,1,ATL 37,0,0,Drew Lock pass complete short right to Daniel Bellinger for 5 yards (tackle by Jessie Bates),2.480,3.450
1,3:37,1,10,ATL 32,0,0,Drew Lock pass complete short left to Wan'Dale Robinson for 9 yards (tackle by Justin Simmons),3.450,4.120
1,2:54,2,1,ATL 23,0,0,Tyrone Tracy left tackle for 5 yards (tackle by Ruke Orhorhoro and Mike Hughes),4.120,4.370
1,2:11,1,10,ATL 18,0,0,Drew Lock pass complete short left to Wan'Dale Robinson for 6 yards (tackle by Lorenzo Carter),4.370,4.810
1,1:30,2,4,ATL 12,0,0,Tyrone Tracy right end for 4 yards (tackle by DeAundre Alford),4.810,5.370
1,0:45,1,8,ATL 8,0,0,Drew Lock pass incomplete short right intended for Wan'Dale Robinson (defended by Jessie Bates),5.370,4.570
1,0:40,2,8,ATL 8,0,0,Darius Slayton right tackle for 6 yards (tackle by DeAundre Alford),4.570,4.950
2,15:00,3,2,ATL 2,6,0,Drew Lock pass complete short left to Tyrone Tracy for 2 yards touchdown,4.950,7.000
2,14:53,,,ATL 15,7,0,Graham Gano kicks extra point good,0.000,0.000
2,14:53,,,NYG 35,7,0,Graham Gano kicks off 65 yards touchback.,0.000,0.940
2,14:53,1,10,ATL 30,7,0,Michael Penix pass complete deep right to Darnell Mooney for 22 yards (tackle by Adoree' Jackson),0.940,2.390
2,14:19,1,10,NYG 48,7,0,Bijan Robinson right tackle for 4 yards (tackle by Raheem Layne),2.390,2.390
2,13:41,2,6,NYG 44,7,0,Tyler Allgeier right tackle for -1 yards (tackle by Boogie Basham),2.390,1.550
2,12:58,3,7,NYG 45,7,0,Michael Penix pass complete short middle to Drake London for 10 yards (tackle by Micah McFadden and Kayvon Thibodeaux),1.550,3.250
2,12:14,1,10,NYG 35,7,0,Michael Penix pass complete short right to Bijan Robinson for -4 yards (tackle by Andru Phillips),3.250,2.160
2,11:32,2,14,NYG 39,7,0,Michael Penix scrambles left guard for 5 yards (tackle by Micah McFadden),2.160,2.150
2,10:46,3,9,NYG 34,7,0,Michael Penix pass incomplete short left intended for Darnell Mooney,2.150,1.060
2,10:41,4,9,NYG 34,7,3,Riley Patterson 52 yard field goal good,1.060,3.000
2,10:36,,,ATL 35,7,3,Bradley Pinion kicks off 65 yards touchback.,0.000,0.940
2,10:36,1,10,NYG 30,7,3,Drew Lock pass incomplete short right intended for Malik Nabers,0.940,0.390
2,10:31,2,10,NYG 30,7,3,Penalty on Evan Neal: False Start 5 yards (accepted) (no play),0.390,-0.280
2,10:31,2,15,NYG 25,7,3,Drew Lock pass complete short right to Jalin Hyatt for 9 yards (tackle by Mike Hughes),-0.280,0.230
2,9:52,3,6,NYG 34,7,3,Drew Lock pass complete short left to Wan'Dale Robinson for 15 yards (tackle by DeAundre Alford and Jessie Bates),0.230,2.190
2,9:06,1,10,NYG 49,7,3,Penalty on Drew Lock: Delay of Game 5 yards (accepted) (no play),2.190,1.860
2,8:51,1,15,NYG 44,7,3,Drew Lock pass complete short right to Wan'Dale Robinson for 8 yards (tackle by AJ Terrell),1.860,2.120
2,8:05,2,6,ATL 48,7,9,Drew Lock pass short left intended for Wan'Dale Robinson is intercepted by Jessie Bates at ATL-45 and returned for 55 yards touchdown,2.120,-7.000
2,7:56,,,NYG 15,7,10,Riley Patterson kicks extra point good,0.000,0.000
2,7:56,,,ATL 35,7,10,Bradley Pinion kicks off 65 yards touchback.,0.000,0.940
2,7:56,1,10,NYG 30,7,10,Tyrone Tracy right tackle for 1 yard (tackle by Kaden Elliss),0.940,0.530
2,7:19,2,9,NYG 31,7,10,Drew Lock pass complete short left to Malik Nabers for 10 yards (tackle by Justin Simmons and Mike Hughes),0.530,1.660
2,6:39,1,10,NYG 41,7,10,Tyrone Tracy left tackle for 3 yards (tackle by Arnold Ebiketie and Eddie Goldman),1.660,1.530
2,6:02,2,7,NYG 44,7,10,Drew Lock sacked by Arnold Ebiketie for -4 yards,1.530,0.300
2,5:20,3,11,NYG 40,7,10,Drew Lock pass incomplete deep middle intended for Malik Nabers,0.300,-0.720
2,5:16,4,11,NYG 40,7,10,Jamie Gillan punts 46 yards fair catch by Avery Williams at ATL-14,-0.720,0.280
2,5:09,1,10,ATL 14,7,10,Michael Penix pass complete short left to Darnell Mooney for 15 yards (tackle by Andru Phillips),-0.280,0.870
2,4:28,1,10,ATL 29,7,10,Bijan Robinson left end for 2 yards (tackle by Rakeem Nunez-Roches and Kayvon Thibodeaux),0.870,0.600
2,3:51,2,8,ATL 31,7,10,Michael Penix pass incomplete short left,0.600,-0.100
2,3:46,3,8,ATL 31,7,10,Michael Penix pass incomplete deep left intended for Darnell Mooney. Penalty on Deonte Banks: Defensive Pass Interference 30 yards (accepted) (no play),-0.100,2.980
2,3:40,1,10,NYG 39,7,10,Tyler Allgeier left tackle for 2 yards (tackle by Darius Muasau and Deonte Banks),2.980,2.710
2,2:58,2,8,NYG 37,7,10,Tyler Allgeier right tackle for 2 yards (tackle by Darius Muasau and Micah McFadden),2.710,2.280
2,2:17,3,6,NYG 35,7,10,Michael Penix pass complete short middle to Darnell Mooney for 19 yards (tackle by Jason Pinnock),2.280,4.510
2,2:00,1,10,NYG 16,7,10,Bijan Robinson right end for 9 yards (tackle by Dane Belton and Tomon Fox),4.510,5.540
2,1:53,,,,,,Timeout #1 by New York Giants,,
2,1:53,2,1,NYG 7,7,10,Bijan Robinson right tackle for 3 yards (tackle by Jordon Riley),5.540,6.280
2,1:48,,,,,,Timeout #2 by New York Giants,,
2,1:48,1,4,NYG 4,7,16,Bijan Robinson left end for 4 yards touchdown,6.280,7.000
2,1:43,,,NYG 15,7,17,Riley Patterson kicks extra point good,0.000,0.000
2,1:43,,,ATL 35,7,17,Bradley Pinion kicks off 61 yards returned by Eric Gray for 37 yards (tackle by DeAngelo Malone and Ross Dwelley),0.000,1.660
2,1:35,1,10,NYG 41,7,17,Drew Lock sacked by Kaden Elliss for -10 yards. Drew Lock fumbles (forced by Kaden Elliss) recovered by Arnold Ebiketie at NYG-31 (tackle by Kaden Elliss),1.660,-3.510
2,1:26,1,10,NYG 31,7,17,Bijan Robinson left end for 3 yards (tackle by Micah McFadden),3.510,3.370
2,1:06,,,,,,Timeout #3 by New York Giants,,
2,1:06,2,7,NYG 28,7,17,Bijan Robinson right end for -1 yards (tackle by Darius Muasau and Cory Durden),3.370,2.540
2,0:30,,,,,,Timeout #1 by Atlanta Falcons,,
2,0:30,3,8,NYG 29,7,17,Michael Penix pass complete short right to Darnell Mooney for 14 yards,2.540,4.580
2,0:27,1,10,NYG 15,7,17,Bijan Robinson right end for -2 yards (tackle by Brian Burns),4.580,3.680
2,0:22,,,,,,Timeout #2 by Atlanta Falcons,,
2,0:22,2,12,NYG 17,7,17,Michael Penix pass complete short right to Drake London for 10 yards (tackle by Raheem Layne),3.680,4.680
2,0:16,,,,,,Timeout #3 by Atlanta Falcons,,
2,0:16,3,2,NYG 7,7,17,Michael Penix pass short right (defended by Dane Belton) intended for Kyle Pitts is intercepted by Cordale Flott in end zone and returned for 26 yards (tackle by Drake London),4.680,-0.610
2,0:07,1,10,NYG 25,7,17,Penalty on Drake London: Personal Foul / Defense 15 yards (accepted) (no play),0.610,1.600
2,0:07,1,10,NYG 40,7,17,Drew Lock pass incomplete short left intended for Daniel Bellinger,1.600,1.050
2,0:04,2,10,NYG 40,7,17,Drew Lock pass incomplete short left intended for Malik Nabers,1.050,0.370
3,15:00,,,ATL 35,7,17,Bradley Pinion kicks off 65 yards touchback.,0.000,0.940
3,15:00,1,10,NYG 30,7,17,Devin Singletary right guard for 3 yards (tackle by David Onyemata),0.940,0.800
3,14:27,2,7,NYG 33,7,23,Drew Lock pass short middle (defended by Zach Harrison) intended for Malik Nabers is intercepted by Matt Judon at NYG-27 and returned for 27 yards touchdown,0.800,-7.000
3,14:20,,,NYG 15,7,24,Riley Patterson kicks extra point good,0.000,0.000
3,14:20,,,ATL 35,7,24,Bradley Pinion kicks off 65 yards touchback.,0.000,0.940
3,14:20,1,10,NYG 30,7,24,Drew Lock pass incomplete short middle,0.940,0.390
3,14:16,2,10,NYG 30,7,24,Tyrone Tracy left tackle for 4 yards (tackle by Zach Harrison and Kaden Elliss),0.390,0.230
3,13:45,3,6,NYG 34,7,24,Drew Lock pass incomplete short right intended for Wan'Dale Robinson (defended by DeAundre Alford),0.230,-1.110
3,13:42,4,6,NYG 34,7,24,Jamie Gillan punts 41 yards returned by Avery Williams for 6 yards (tackle by Dane Belton and Casey Kreiter),-1.110,-1.000
3,13:31,1,10,ATL 31,7,24,Bijan Robinson right guard for 14 yards (tackle by Jason Pinnock and Dane Belton),1.000,1.930
3,12:50,1,10,ATL 45,7,24,Bijan Robinson right end for -1 yards (tackle by Ty Summers),1.930,1.250
3,12:13,2,11,ATL 44,7,24,Michael Penix pass complete short middle to Drake London for 15 yards (tackle by Raheem Layne),1.250,2.850
3,11:26,1,10,NYG 41,7,24,Tyler Allgeier left end for 12 yards (tackle by Deonte Banks),2.850,3.640
3,10:43,1,10,NYG 29,7,24,Michael Penix pass incomplete short left intended for Charlie Woerner,3.640,3.100
3,10:37,2,10,NYG 29,7,24,Michael Penix pass complete short left to Tyler Allgeier for 9 yards (tackle by Ty Summers),3.100,3.600
3,10:08,3,1,NYG 20,7,24,Tyler Allgeier left tackle for 2 yards (tackle by Cory Durden and Boogie Basham),3.600,4.370
3,9:31,1,10,NYG 18,7,24,Bijan Robinson right tackle for 3 yards (tackle by Cory Durden),4.370,4.250
3,8:50,2,7,NYG 15,7,24,Bijan Robinson right guard for no gain (tackle by Andru Phillips and Boogie Basham),4.250,3.580
3,8:08,3,6,NYG 15,7,24,Michael Penix pass complete short right to Bijan Robinson for 13 yards (tackle by Ty Summers),3.580,6.740
3,7:23,1,2,NYG 2,7,24,Michael Penix pass incomplete short left intended for Drake London (defended by Deonte Banks),6.740,5.720
3,7:19,2,2,NYG 2,7,30,Bijan Robinson left end for 2 yards touchdown,5.720,7.000
3,7:14,,,NYG 15,7,31,Riley Patterson kicks extra point good,0.000,0.000
3,7:14,,,ATL 35,7,31,Bradley Pinion kicks off 65 yards touchback.,0.000,0.940
3,7:14,1,10,NYG 30,7,31,Drew Lock pass complete short right to Malik Nabers for 6 yards (tackle by DeAundre Alford),0.940,1.200
3,6:41,2,4,NYG 36,7,31,Devin Singletary right tackle for no gain (tackle by Zach Harrison and Kaden Elliss),1.200,0.500
3,6:02,3,4,NYG 36,7,31,Drew Lock pass incomplete short left intended for Wan'Dale Robinson (defended by DeAundre Alford),0.500,-0.980
3,5:58,4,4,NYG 36,7,31,Jamie Gillan punts 51 yards fair catch by Avery Williams at ATL-13,-0.980,0.320
3,5:51,1,10,ATL 13,7,31,Tyler Allgeier left end for 2 yards (tackle by Darius Muasau and Tomon Fox),-0.320,-0.570
3,5:13,2,8,ATL 15,7,31,Michael Penix pass complete short right to Ray-Ray McCloud for 7 yards (tackle by Darius Muasau),-0.570,-0.350
3,4:30,3,1,ATL 22,7,31,Tyler Allgeier left guard for 1 yard (tackle by Cory Durden and Andru Phillips),-0.350,0.480
3,3:51,1,10,ATL 23,7,31,Tyler Allgeier left end for 4 yards (tackle by Darius Muasau),0.480,0.470
3,3:09,2,6,ATL 27,7,31,Michael Penix pass complete short middle to Ray-Ray McCloud for 8 yards (tackle by Cordale Flott),0.470,1.270
3,2:30,1,10,ATL 35,7,31,Bijan Robinson right tackle for 1 yard (tackle by Ty Summers and Cory Durden),1.270,0.860
3,1:49,2,9,ATL 36,7,31,Bijan Robinson right tackle for 11 yards (tackle by Dane Belton and Ty Summers),0.860,2.060
3,1:06,1,10,ATL 47,7,31,Michael Penix pass complete deep middle to Chris Blair for 17 yards (tackle by Jason Pinnock),2.060,3.180
3,0:22,1,10,NYG 36,7,31,Bijan Robinson left tackle for 8 yards (tackle by Dane Belton),3.180,3.720
4,15:00,2,2,NYG 28,7,31,Bijan Robinson left tackle for 1 yard (tackle by Darius Muasau and Ty Summers),3.720,3.140
4,14:16,3,1,NYG 27,7,31,Bijan Robinson left tackle for 6 yards (tackle by Jason Pinnock),3.140,4.170
4,13:32,1,10,NYG 21,7,31,Tyler Allgeier left end for 2 yards (tackle by Brian Burns),4.170,3.900
4,12:48,2,8,NYG 19,7,31,Michael Penix pass complete short right to Kyle Pitts for 7 yards (tackle by Jason Pinnock and Darius Muasau),3.900,4.490
4,12:03,3,1,NYG 12,7,31,Bijan Robinson left end for no gain (tackle by Cordale Flott). Penalty on Drew Dalman: Offensive Holding 10 yards (accepted) (no play),4.490,2.810
4,11:32,3,11,NYG 22,7,31,Michael Penix pass complete short right to Ray-Ray McCloud for 4 yards (tackle by Cordale Flott),2.810,2.250
4,10:50,4,7,NYG 18,7,34,Riley Patterson 37 yard field goal good,2.250,3.000
4,10:47,,,ATL 35,7,34,Bradley Pinion kicks off 65 yards touchback.,0.000,0.940
4,10:47,1,10,NYG 30,7,34,Drew Lock pass incomplete short right intended for Malik Nabers (defended by Mike Hughes),0.940,0.390
4,10:41,2,10,NYG 30,7,34,Drew Lock pass complete short right to Tyrone Tracy for 16 yards (tackle by Arnold Ebiketie),0.390,1.990
4,9:58,1,10,NYG 46,7,34,Drew Lock pass incomplete deep right intended for Jalin Hyatt,1.990,1.450
4,9:53,2,10,NYG 46,7,34,Drew Lock right tackle for 1 yard (tackle by Arnold Ebiketie and Grady Jarrett),1.450,0.890
4,9:09,3,9,NYG 47,7,34,Penalty on Matt Judon: Defensive Offside 5 yards (accepted) (no play),0.890,1.550
4,8:44,3,4,ATL 48,7,34,Drew Lock pass complete deep right to Malik Nabers for no gain. Penalty on Malik Nabers: Illegal Shift 5 yards (accepted) (no play),1.550,0.890
4,8:16,3,9,NYG 47,7,34,Drew Lock sacked by Matt Judon for -7 yards,0.890,-0.720
4,7:32,4,16,NYG 40,7,34,Jamie Gillan punts 21 yards downed by Ty Summers,-0.720,-1.530
4,7:23,1,10,ATL 39,7,34,Tyler Allgeier left tackle for -3 yards (tackle by Jason Pinnock and Ty Summers). Penalty on Matthew Bergeron: Offensive Holding 10 yards (declined),1.530,0.580
4,7:01,2,13,ATL 36,7,34,Tyler Allgeier left end for -1 yards (tackle by Elijah Garcia and Andru Phillips),0.580,-0.230
4,6:14,3,14,ATL 35,7,34,Michael Penix pass complete short right to Darnell Mooney for 12 yards (tackle by Cordale Flott),-0.230,-0.260
4,5:32,4,2,ATL 47,7,34,Bradley Pinion punts 42 yards fair catch by Ihmir Smith-Marsette at NYG-11,-0.260,0.370
4,5:26,1,10,NYG 11,7,34,Drew Lock pass complete short right to Malik Nabers for 5 yards (tackle by JD Bertrand),-0.370,-0.300
4,4:51,2,5,NYG 16,7,34,Drew Lock pass complete short left to Wan'Dale Robinson for 9 yards (tackle by JD Bertrand),-0.300,0.610
4,4:23,1,10,NYG 25,7,34,Drew Lock pass complete short left to Darius Slayton for 21 yards (tackle by JD Bertrand),0.610,1.990
4,4:13,1,10,NYG 46,7,34,Drew Lock pass complete short right to Wan'Dale Robinson for 11 yards (tackle by JD Bertrand and Nathan Landman),1.990,2.720
4,3:42,1,10,ATL 43,7,34,Drew Lock pass complete short left to Eric Gray for 2 yards (tackle by Kevin King),2.720,2.450
4,3:22,2,8,ATL 41,7,34,Drew Lock pass complete short left to Tyrone Tracy for 16 yards (tackle by Nathan Landman and Arnold Ebiketie),2.450,3.910
4,2:45,1,10,ATL 25,7,34,Penalty on Jermaine Eluemunor: False Start 5 yards (accepted) (no play),3.910,3.580
4,2:45,1,15,ATL 30,7,34,Drew Lock pass complete short left to Malik Nabers for no gain (tackle by Mike Hughes). Penalty on John Michael Schmitz: Offensive Holding 10 yards (accepted) (no play),3.580,2.920
4,2:40,1,25,ATL 40,7,34,Drew Lock pass complete short left to Malik Nabers for 14 yards (tackle by Nathan Landman and Mike Hughes),2.920,3.230
4,2:10,2,11,ATL 26,7,34,Drew Lock pass complete deep left to Malik Nabers for 21 yards (tackle by Mike Hughes). Penalty on Natrone Brooks: Defensive Offside 5 yards (declined),3.230,6.060
4,2:04,1,5,ATL 5,7,34,Tyrone Tracy right end for no gain touchdown. Penalty on Wan'Dale Robinson: Offensive Holding 10 yards (accepted) (no play),6.060,4.370
4,1:59,1,15,ATL 15,7,34,Drew Lock pass complete short right to Wan'Dale Robinson for 4 yards (tackle by Kentavius Street and Nathan Landman),4.370,4.020
4,1:33,2,11,ATL 11,7,34,Penalty on Evan Neal: False Start 5 yards (accepted) (no play),4.020,3.340
4,1:33,,,,,,Timeout #1 by New York Giants,,
4,1:33,2,16,ATL 16,7,34,Drew Lock pass incomplete deep left intended for Malik Nabers (defended by Mike Hughes),3.340,2.850
4,1:28,3,16,ATL 16,7,34,Drew Lock pass incomplete deep right intended for Malik Nabers (defended by Clark Phillips),2.850,2.380
4,1:22,,,,,,Timeout #1 by Atlanta Falcons,,
4,1:22,4,16,ATL 16,7,34,Penalty on Evan Neal: False Start 5 yards (accepted) (no play),2.380,2.060
4,1:22,4,21,ATL 21,7,34,Drew Lock pass incomplete deep right intended for Darius Slayton,2.060,-0.410
4,1:12,1,10,ATL 22,7,34,Michael Penix kneels for -1 yards,0.410,-0.270
4,0:31,2,11,ATL 21,7,34,Michael Penix kneels for -2 yards,-0.270,-1.290